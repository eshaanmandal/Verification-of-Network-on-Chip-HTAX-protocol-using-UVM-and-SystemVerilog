///////////////////////////////////////////////////////////////////////////
// Texas A&M University
// CSCE 616 Hardware Design Verification
// Created by  : Prof. Quinn and Saumil Gogri
///////////////////////////////////////////////////////////////////////////

`include "base_test.sv"
`include "simple_random_test.sv"
`include "multiport_sequential_random_test.sv"
`include "multiport_parallel_random_test.sv"
`include "variable_delay_test.sv"
`include "packet_length_test.sv"
